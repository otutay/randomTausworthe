-------------------------------------------------------------------------------
-- Title      : Noise packge
-- Project    : noise generator
-------------------------------------------------------------------------------
-- File       : noisePckg.vhd
-- Author     : osmant  <otutaysalgir@gmail.com>
-- Company    :
-- Created    : 2019-09-08
-- Last update: 2019-09-08
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------
-- Copyright (c) 2019
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-09-08  1.0      osmant  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package noisePackage is
  constant c_dataBitW : integer := 32;


end package noisePackage;

package body noisePackage is

end package body noisePackage;
